module transmitter(
    input wire clk,
    input wire [7:0] data,
    input wire is_addr,
    input wire send_en,
    output wire sda,
    output wire scl
);

endmodule