module imu_data_acquisition(input clk);

    always @(posedge clk) begin

    end

endmodule